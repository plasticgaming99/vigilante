module main

import time

fn main() {
	time.sleep(1*time.second)
}