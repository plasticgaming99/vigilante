module quickev
