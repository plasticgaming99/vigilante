// quickev is a single threaded event loop librrary
// not recommended for using in network applications

module quickev
