module main

// logger???
// like [  OK  ]?
// [*     ]
// [**    ]
// [ ***  ]
// [  *** ]
// [   ***]
// [    **]
// [     *]
// [FAILED]
